module tb_ajw_addsub_unit;
    // TODO: Create TB to verify our CLA.......
endmodule
